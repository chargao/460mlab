module KeyboardController (PS2CLK,DATA);
input PS2CLK;
input DATA;


endmodule
